`include "include.vh"

/*
--------------------------------
module reg_manage
・レジスタを管理
・データハザードの検出
--------------------------------
*/
