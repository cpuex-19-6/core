`include "include.vh"

`default_nettype none

module uart_input_generate #(
    CLK_FREQ = `CLK_PER_SEC, BAUD = `DEFAULT_BAUD)(
        output wire rx,
        input  wire clk,
        input  wire rstn);

    wire [8-1:0] to_send[1300-1:0];
    assign to_send[0] = 8'hc2;
    assign to_send[1] = 8'h8c;
    assign to_send[2] = 8'h00;
    assign to_send[3] = 8'h00;
    assign to_send[4] = 8'h42;
    assign to_send[5] = 8'h0c;
    assign to_send[6] = 8'h00;
    assign to_send[7] = 8'h00;
    assign to_send[8] = 8'hc1;
    assign to_send[9] = 8'ha0;
    assign to_send[10] = 8'h00;
    assign to_send[11] = 8'h00;
    assign to_send[12] = 8'h41;
    assign to_send[13] = 8'ha0;
    assign to_send[14] = 8'h00;
    assign to_send[15] = 8'h00;
    assign to_send[16] = 8'h41;
    assign to_send[17] = 8'hf0;
    assign to_send[18] = 8'h00;
    assign to_send[19] = 8'h00;
    assign to_send[20] = 8'h3f;
    assign to_send[21] = 8'h80;
    assign to_send[22] = 8'h00;
    assign to_send[23] = 8'h00;
    assign to_send[24] = 8'h42;
    assign to_send[25] = 8'h48;
    assign to_send[26] = 8'h00;
    assign to_send[27] = 8'h00;
    assign to_send[28] = 8'h42;
    assign to_send[29] = 8'h48;
    assign to_send[30] = 8'h00;
    assign to_send[31] = 8'h00;
    assign to_send[32] = 8'h43;
    assign to_send[33] = 8'h7f;
    assign to_send[34] = 8'h00;
    assign to_send[35] = 8'h00;
    assign to_send[36] = 8'h00;
    assign to_send[37] = 8'h00;
    assign to_send[38] = 8'h00;
    assign to_send[39] = 8'h00;
    assign to_send[40] = 8'h00;
    assign to_send[41] = 8'h00;
    assign to_send[42] = 8'h00;
    assign to_send[43] = 8'h01;
    assign to_send[44] = 8'h00;
    assign to_send[45] = 8'h00;
    assign to_send[46] = 8'h00;
    assign to_send[47] = 8'h01;
    assign to_send[48] = 8'h00;
    assign to_send[49] = 8'h00;
    assign to_send[50] = 8'h00;
    assign to_send[51] = 8'h00;
    assign to_send[52] = 8'h41;
    assign to_send[53] = 8'ha0;
    assign to_send[54] = 8'h00;
    assign to_send[55] = 8'h00;
    assign to_send[56] = 8'h41;
    assign to_send[57] = 8'ha0;
    assign to_send[58] = 8'h00;
    assign to_send[59] = 8'h00;
    assign to_send[60] = 8'h42;
    assign to_send[61] = 8'h82;
    assign to_send[62] = 8'h00;
    assign to_send[63] = 8'h00;
    assign to_send[64] = 8'h00;
    assign to_send[65] = 8'h00;
    assign to_send[66] = 8'h00;
    assign to_send[67] = 8'h00;
    assign to_send[68] = 8'h41;
    assign to_send[69] = 8'ha0;
    assign to_send[70] = 8'h00;
    assign to_send[71] = 8'h00;
    assign to_send[72] = 8'h42;
    assign to_send[73] = 8'h34;
    assign to_send[74] = 8'h00;
    assign to_send[75] = 8'h00;
    assign to_send[76] = 8'h3f;
    assign to_send[77] = 8'h80;
    assign to_send[78] = 8'h00;
    assign to_send[79] = 8'h00;
    assign to_send[80] = 8'h3f;
    assign to_send[81] = 8'h80;
    assign to_send[82] = 8'h00;
    assign to_send[83] = 8'h00;
    assign to_send[84] = 8'h43;
    assign to_send[85] = 8'h7a;
    assign to_send[86] = 8'h00;
    assign to_send[87] = 8'h00;
    assign to_send[88] = 8'h43;
    assign to_send[89] = 8'h00;
    assign to_send[90] = 8'h00;
    assign to_send[91] = 8'h00;
    assign to_send[92] = 8'h43;
    assign to_send[93] = 8'h52;
    assign to_send[94] = 8'h00;
    assign to_send[95] = 8'h00;
    assign to_send[96] = 8'h00;
    assign to_send[97] = 8'h00;
    assign to_send[98] = 8'h00;
    assign to_send[99] = 8'h00;
    assign to_send[100] = 8'h00;
    assign to_send[101] = 8'h00;
    assign to_send[102] = 8'h00;
    assign to_send[103] = 8'h00;
    assign to_send[104] = 8'h00;
    assign to_send[105] = 8'h00;
    assign to_send[106] = 8'h00;
    assign to_send[107] = 8'h03;
    assign to_send[108] = 8'h00;
    assign to_send[109] = 8'h00;
    assign to_send[110] = 8'h00;
    assign to_send[111] = 8'h01;
    assign to_send[112] = 8'h00;
    assign to_send[113] = 8'h00;
    assign to_send[114] = 8'h00;
    assign to_send[115] = 8'h00;
    assign to_send[116] = 8'h41;
    assign to_send[117] = 8'hc8;
    assign to_send[118] = 8'h00;
    assign to_send[119] = 8'h00;
    assign to_send[120] = 8'h42;
    assign to_send[121] = 8'h20;
    assign to_send[122] = 8'h00;
    assign to_send[123] = 8'h00;
    assign to_send[124] = 8'h42;
    assign to_send[125] = 8'h8c;
    assign to_send[126] = 8'h00;
    assign to_send[127] = 8'h00;
    assign to_send[128] = 8'h00;
    assign to_send[129] = 8'h00;
    assign to_send[130] = 8'h00;
    assign to_send[131] = 8'h00;
    assign to_send[132] = 8'h00;
    assign to_send[133] = 8'h00;
    assign to_send[134] = 8'h00;
    assign to_send[135] = 8'h00;
    assign to_send[136] = 8'h42;
    assign to_send[137] = 8'h20;
    assign to_send[138] = 8'h00;
    assign to_send[139] = 8'h00;
    assign to_send[140] = 8'h3f;
    assign to_send[141] = 8'h80;
    assign to_send[142] = 8'h00;
    assign to_send[143] = 8'h00;
    assign to_send[144] = 8'h3f;
    assign to_send[145] = 8'h80;
    assign to_send[146] = 8'h00;
    assign to_send[147] = 8'h00;
    assign to_send[148] = 8'h43;
    assign to_send[149] = 8'h7a;
    assign to_send[150] = 8'h00;
    assign to_send[151] = 8'h00;
    assign to_send[152] = 8'h43;
    assign to_send[153] = 8'h00;
    assign to_send[154] = 8'h00;
    assign to_send[155] = 8'h00;
    assign to_send[156] = 8'h43;
    assign to_send[157] = 8'h52;
    assign to_send[158] = 8'h00;
    assign to_send[159] = 8'h00;
    assign to_send[160] = 8'h00;
    assign to_send[161] = 8'h00;
    assign to_send[162] = 8'h00;
    assign to_send[163] = 8'h00;
    assign to_send[164] = 8'h00;
    assign to_send[165] = 8'h00;
    assign to_send[166] = 8'h00;
    assign to_send[167] = 8'h00;
    assign to_send[168] = 8'h00;
    assign to_send[169] = 8'h00;
    assign to_send[170] = 8'h00;
    assign to_send[171] = 8'h03;
    assign to_send[172] = 8'h00;
    assign to_send[173] = 8'h00;
    assign to_send[174] = 8'h00;
    assign to_send[175] = 8'h01;
    assign to_send[176] = 8'h00;
    assign to_send[177] = 8'h00;
    assign to_send[178] = 8'h00;
    assign to_send[179] = 8'h00;
    assign to_send[180] = 8'h00;
    assign to_send[181] = 8'h00;
    assign to_send[182] = 8'h00;
    assign to_send[183] = 8'h00;
    assign to_send[184] = 8'h41;
    assign to_send[185] = 8'hf0;
    assign to_send[186] = 8'h00;
    assign to_send[187] = 8'h00;
    assign to_send[188] = 8'h41;
    assign to_send[189] = 8'hf0;
    assign to_send[190] = 8'h00;
    assign to_send[191] = 8'h00;
    assign to_send[192] = 8'h00;
    assign to_send[193] = 8'h00;
    assign to_send[194] = 8'h00;
    assign to_send[195] = 8'h00;
    assign to_send[196] = 8'hc0;
    assign to_send[197] = 8'ha0;
    assign to_send[198] = 8'h00;
    assign to_send[199] = 8'h00;
    assign to_send[200] = 8'h00;
    assign to_send[201] = 8'h00;
    assign to_send[202] = 8'h00;
    assign to_send[203] = 8'h00;
    assign to_send[204] = 8'hbf;
    assign to_send[205] = 8'h80;
    assign to_send[206] = 8'h00;
    assign to_send[207] = 8'h00;
    assign to_send[208] = 8'h3f;
    assign to_send[209] = 8'h80;
    assign to_send[210] = 8'h00;
    assign to_send[211] = 8'h00;
    assign to_send[212] = 8'h43;
    assign to_send[213] = 8'h7a;
    assign to_send[214] = 8'h00;
    assign to_send[215] = 8'h00;
    assign to_send[216] = 8'h43;
    assign to_send[217] = 8'h00;
    assign to_send[218] = 8'h00;
    assign to_send[219] = 8'h00;
    assign to_send[220] = 8'h43;
    assign to_send[221] = 8'h53;
    assign to_send[222] = 8'h00;
    assign to_send[223] = 8'h00;
    assign to_send[224] = 8'h00;
    assign to_send[225] = 8'h00;
    assign to_send[226] = 8'h00;
    assign to_send[227] = 8'h00;
    assign to_send[228] = 8'h00;
    assign to_send[229] = 8'h00;
    assign to_send[230] = 8'h00;
    assign to_send[231] = 8'h00;
    assign to_send[232] = 8'h00;
    assign to_send[233] = 8'h00;
    assign to_send[234] = 8'h00;
    assign to_send[235] = 8'h01;
    assign to_send[236] = 8'h00;
    assign to_send[237] = 8'h00;
    assign to_send[238] = 8'h00;
    assign to_send[239] = 8'h01;
    assign to_send[240] = 8'h00;
    assign to_send[241] = 8'h00;
    assign to_send[242] = 8'h00;
    assign to_send[243] = 8'h00;
    assign to_send[244] = 8'h41;
    assign to_send[245] = 8'ha0;
    assign to_send[246] = 8'h00;
    assign to_send[247] = 8'h00;
    assign to_send[248] = 8'h41;
    assign to_send[249] = 8'h20;
    assign to_send[250] = 8'h00;
    assign to_send[251] = 8'h00;
    assign to_send[252] = 8'h41;
    assign to_send[253] = 8'hf0;
    assign to_send[254] = 8'h00;
    assign to_send[255] = 8'h00;
    assign to_send[256] = 8'h00;
    assign to_send[257] = 8'h00;
    assign to_send[258] = 8'h00;
    assign to_send[259] = 8'h00;
    assign to_send[260] = 8'hc1;
    assign to_send[261] = 8'h20;
    assign to_send[262] = 8'h00;
    assign to_send[263] = 8'h00;
    assign to_send[264] = 8'h42;
    assign to_send[265] = 8'ha0;
    assign to_send[266] = 8'h00;
    assign to_send[267] = 8'h00;
    assign to_send[268] = 8'h3f;
    assign to_send[269] = 8'h80;
    assign to_send[270] = 8'h00;
    assign to_send[271] = 8'h00;
    assign to_send[272] = 8'h3f;
    assign to_send[273] = 8'h80;
    assign to_send[274] = 8'h00;
    assign to_send[275] = 8'h00;
    assign to_send[276] = 8'h43;
    assign to_send[277] = 8'h7a;
    assign to_send[278] = 8'h00;
    assign to_send[279] = 8'h00;
    assign to_send[280] = 8'h43;
    assign to_send[281] = 8'h00;
    assign to_send[282] = 8'h00;
    assign to_send[283] = 8'h00;
    assign to_send[284] = 8'h43;
    assign to_send[285] = 8'h53;
    assign to_send[286] = 8'h00;
    assign to_send[287] = 8'h00;
    assign to_send[288] = 8'h00;
    assign to_send[289] = 8'h00;
    assign to_send[290] = 8'h00;
    assign to_send[291] = 8'h00;
    assign to_send[292] = 8'h00;
    assign to_send[293] = 8'h00;
    assign to_send[294] = 8'h00;
    assign to_send[295] = 8'h00;
    assign to_send[296] = 8'h00;
    assign to_send[297] = 8'h00;
    assign to_send[298] = 8'h00;
    assign to_send[299] = 8'h02;
    assign to_send[300] = 8'h00;
    assign to_send[301] = 8'h00;
    assign to_send[302] = 8'h00;
    assign to_send[303] = 8'h01;
    assign to_send[304] = 8'h00;
    assign to_send[305] = 8'h00;
    assign to_send[306] = 8'h00;
    assign to_send[307] = 8'h00;
    assign to_send[308] = 8'h00;
    assign to_send[309] = 8'h00;
    assign to_send[310] = 8'h00;
    assign to_send[311] = 8'h00;
    assign to_send[312] = 8'hbf;
    assign to_send[313] = 8'hc0;
    assign to_send[314] = 8'h00;
    assign to_send[315] = 8'h00;
    assign to_send[316] = 8'hbf;
    assign to_send[317] = 8'h80;
    assign to_send[318] = 8'h00;
    assign to_send[319] = 8'h00;
    assign to_send[320] = 8'h00;
    assign to_send[321] = 8'h00;
    assign to_send[322] = 8'h00;
    assign to_send[323] = 8'h00;
    assign to_send[324] = 8'h00;
    assign to_send[325] = 8'h00;
    assign to_send[326] = 8'h00;
    assign to_send[327] = 8'h00;
    assign to_send[328] = 8'h42;
    assign to_send[329] = 8'h48;
    assign to_send[330] = 8'h00;
    assign to_send[331] = 8'h00;
    assign to_send[332] = 8'h3f;
    assign to_send[333] = 8'h80;
    assign to_send[334] = 8'h00;
    assign to_send[335] = 8'h00;
    assign to_send[336] = 8'h3f;
    assign to_send[337] = 8'h80;
    assign to_send[338] = 8'h00;
    assign to_send[339] = 8'h00;
    assign to_send[340] = 8'h43;
    assign to_send[341] = 8'h7a;
    assign to_send[342] = 8'h00;
    assign to_send[343] = 8'h00;
    assign to_send[344] = 8'h43;
    assign to_send[345] = 8'h00;
    assign to_send[346] = 8'h00;
    assign to_send[347] = 8'h00;
    assign to_send[348] = 8'h43;
    assign to_send[349] = 8'h53;
    assign to_send[350] = 8'h00;
    assign to_send[351] = 8'h00;
    assign to_send[352] = 8'h00;
    assign to_send[353] = 8'h00;
    assign to_send[354] = 8'h00;
    assign to_send[355] = 8'h00;
    assign to_send[356] = 8'h00;
    assign to_send[357] = 8'h00;
    assign to_send[358] = 8'h00;
    assign to_send[359] = 8'h00;
    assign to_send[360] = 8'h00;
    assign to_send[361] = 8'h00;
    assign to_send[362] = 8'h00;
    assign to_send[363] = 8'h01;
    assign to_send[364] = 8'h00;
    assign to_send[365] = 8'h00;
    assign to_send[366] = 8'h00;
    assign to_send[367] = 8'h01;
    assign to_send[368] = 8'h00;
    assign to_send[369] = 8'h00;
    assign to_send[370] = 8'h00;
    assign to_send[371] = 8'h00;
    assign to_send[372] = 8'h41;
    assign to_send[373] = 8'hb0;
    assign to_send[374] = 8'h00;
    assign to_send[375] = 8'h00;
    assign to_send[376] = 8'h41;
    assign to_send[377] = 8'he0;
    assign to_send[378] = 8'h00;
    assign to_send[379] = 8'h00;
    assign to_send[380] = 8'h41;
    assign to_send[381] = 8'he0;
    assign to_send[382] = 8'h00;
    assign to_send[383] = 8'h00;
    assign to_send[384] = 8'h00;
    assign to_send[385] = 8'h00;
    assign to_send[386] = 8'h00;
    assign to_send[387] = 8'h00;
    assign to_send[388] = 8'hc0;
    assign to_send[389] = 8'ha0;
    assign to_send[390] = 8'h00;
    assign to_send[391] = 8'h00;
    assign to_send[392] = 8'h00;
    assign to_send[393] = 8'h00;
    assign to_send[394] = 8'h00;
    assign to_send[395] = 8'h00;
    assign to_send[396] = 8'h3f;
    assign to_send[397] = 8'h80;
    assign to_send[398] = 8'h00;
    assign to_send[399] = 8'h00;
    assign to_send[400] = 8'h3f;
    assign to_send[401] = 8'h80;
    assign to_send[402] = 8'h00;
    assign to_send[403] = 8'h00;
    assign to_send[404] = 8'h43;
    assign to_send[405] = 8'h7a;
    assign to_send[406] = 8'h00;
    assign to_send[407] = 8'h00;
    assign to_send[408] = 8'h00;
    assign to_send[409] = 8'h00;
    assign to_send[410] = 8'h00;
    assign to_send[411] = 8'h00;
    assign to_send[412] = 8'h43;
    assign to_send[413] = 8'h53;
    assign to_send[414] = 8'h00;
    assign to_send[415] = 8'h00;
    assign to_send[416] = 8'h43;
    assign to_send[417] = 8'h53;
    assign to_send[418] = 8'h00;
    assign to_send[419] = 8'h00;
    assign to_send[420] = 8'h00;
    assign to_send[421] = 8'h00;
    assign to_send[422] = 8'h00;
    assign to_send[423] = 8'h00;
    assign to_send[424] = 8'h00;
    assign to_send[425] = 8'h00;
    assign to_send[426] = 8'h00;
    assign to_send[427] = 8'h03;
    assign to_send[428] = 8'h00;
    assign to_send[429] = 8'h00;
    assign to_send[430] = 8'h00;
    assign to_send[431] = 8'h01;
    assign to_send[432] = 8'h00;
    assign to_send[433] = 8'h00;
    assign to_send[434] = 8'h00;
    assign to_send[435] = 8'h00;
    assign to_send[436] = 8'h42;
    assign to_send[437] = 8'h20;
    assign to_send[438] = 8'h00;
    assign to_send[439] = 8'h00;
    assign to_send[440] = 8'h41;
    assign to_send[441] = 8'he0;
    assign to_send[442] = 8'h00;
    assign to_send[443] = 8'h00;
    assign to_send[444] = 8'h41;
    assign to_send[445] = 8'he0;
    assign to_send[446] = 8'h00;
    assign to_send[447] = 8'h00;
    assign to_send[448] = 8'h00;
    assign to_send[449] = 8'h00;
    assign to_send[450] = 8'h00;
    assign to_send[451] = 8'h00;
    assign to_send[452] = 8'hc0;
    assign to_send[453] = 8'ha0;
    assign to_send[454] = 8'h00;
    assign to_send[455] = 8'h00;
    assign to_send[456] = 8'h00;
    assign to_send[457] = 8'h00;
    assign to_send[458] = 8'h00;
    assign to_send[459] = 8'h00;
    assign to_send[460] = 8'h3f;
    assign to_send[461] = 8'h80;
    assign to_send[462] = 8'h00;
    assign to_send[463] = 8'h00;
    assign to_send[464] = 8'h3f;
    assign to_send[465] = 8'h80;
    assign to_send[466] = 8'h00;
    assign to_send[467] = 8'h00;
    assign to_send[468] = 8'h43;
    assign to_send[469] = 8'h7a;
    assign to_send[470] = 8'h00;
    assign to_send[471] = 8'h00;
    assign to_send[472] = 8'h00;
    assign to_send[473] = 8'h00;
    assign to_send[474] = 8'h00;
    assign to_send[475] = 8'h00;
    assign to_send[476] = 8'h43;
    assign to_send[477] = 8'h53;
    assign to_send[478] = 8'h00;
    assign to_send[479] = 8'h00;
    assign to_send[480] = 8'h43;
    assign to_send[481] = 8'h53;
    assign to_send[482] = 8'h00;
    assign to_send[483] = 8'h00;
    assign to_send[484] = 8'h00;
    assign to_send[485] = 8'h00;
    assign to_send[486] = 8'h00;
    assign to_send[487] = 8'h00;
    assign to_send[488] = 8'h00;
    assign to_send[489] = 8'h00;
    assign to_send[490] = 8'h00;
    assign to_send[491] = 8'h03;
    assign to_send[492] = 8'h00;
    assign to_send[493] = 8'h00;
    assign to_send[494] = 8'h00;
    assign to_send[495] = 8'h01;
    assign to_send[496] = 8'h00;
    assign to_send[497] = 8'h00;
    assign to_send[498] = 8'h00;
    assign to_send[499] = 8'h00;
    assign to_send[500] = 8'h00;
    assign to_send[501] = 8'h00;
    assign to_send[502] = 8'h00;
    assign to_send[503] = 8'h00;
    assign to_send[504] = 8'h41;
    assign to_send[505] = 8'h70;
    assign to_send[506] = 8'h00;
    assign to_send[507] = 8'h00;
    assign to_send[508] = 8'h41;
    assign to_send[509] = 8'h70;
    assign to_send[510] = 8'h00;
    assign to_send[511] = 8'h00;
    assign to_send[512] = 8'h00;
    assign to_send[513] = 8'h00;
    assign to_send[514] = 8'h00;
    assign to_send[515] = 8'h00;
    assign to_send[516] = 8'hc0;
    assign to_send[517] = 8'ha0;
    assign to_send[518] = 8'h00;
    assign to_send[519] = 8'h00;
    assign to_send[520] = 8'h00;
    assign to_send[521] = 8'h00;
    assign to_send[522] = 8'h00;
    assign to_send[523] = 8'h00;
    assign to_send[524] = 8'hbf;
    assign to_send[525] = 8'h80;
    assign to_send[526] = 8'h00;
    assign to_send[527] = 8'h00;
    assign to_send[528] = 8'h3f;
    assign to_send[529] = 8'h80;
    assign to_send[530] = 8'h00;
    assign to_send[531] = 8'h00;
    assign to_send[532] = 8'h43;
    assign to_send[533] = 8'h7a;
    assign to_send[534] = 8'h00;
    assign to_send[535] = 8'h00;
    assign to_send[536] = 8'h00;
    assign to_send[537] = 8'h00;
    assign to_send[538] = 8'h00;
    assign to_send[539] = 8'h00;
    assign to_send[540] = 8'h43;
    assign to_send[541] = 8'h53;
    assign to_send[542] = 8'h00;
    assign to_send[543] = 8'h00;
    assign to_send[544] = 8'h43;
    assign to_send[545] = 8'h53;
    assign to_send[546] = 8'h00;
    assign to_send[547] = 8'h00;
    assign to_send[548] = 8'h00;
    assign to_send[549] = 8'h00;
    assign to_send[550] = 8'h00;
    assign to_send[551] = 8'h00;
    assign to_send[552] = 8'h00;
    assign to_send[553] = 8'h00;
    assign to_send[554] = 8'h00;
    assign to_send[555] = 8'h03;
    assign to_send[556] = 8'h00;
    assign to_send[557] = 8'h00;
    assign to_send[558] = 8'h00;
    assign to_send[559] = 8'h01;
    assign to_send[560] = 8'h00;
    assign to_send[561] = 8'h00;
    assign to_send[562] = 8'h00;
    assign to_send[563] = 8'h00;
    assign to_send[564] = 8'h41;
    assign to_send[565] = 8'h70;
    assign to_send[566] = 8'h00;
    assign to_send[567] = 8'h00;
    assign to_send[568] = 8'h41;
    assign to_send[569] = 8'hc8;
    assign to_send[570] = 8'h00;
    assign to_send[571] = 8'h00;
    assign to_send[572] = 8'h41;
    assign to_send[573] = 8'hc8;
    assign to_send[574] = 8'h00;
    assign to_send[575] = 8'h00;
    assign to_send[576] = 8'h00;
    assign to_send[577] = 8'h00;
    assign to_send[578] = 8'h00;
    assign to_send[579] = 8'h00;
    assign to_send[580] = 8'hc0;
    assign to_send[581] = 8'ha0;
    assign to_send[582] = 8'h00;
    assign to_send[583] = 8'h00;
    assign to_send[584] = 8'h42;
    assign to_send[585] = 8'h8c;
    assign to_send[586] = 8'h00;
    assign to_send[587] = 8'h00;
    assign to_send[588] = 8'h3f;
    assign to_send[589] = 8'h80;
    assign to_send[590] = 8'h00;
    assign to_send[591] = 8'h00;
    assign to_send[592] = 8'h3f;
    assign to_send[593] = 8'h80;
    assign to_send[594] = 8'h00;
    assign to_send[595] = 8'h00;
    assign to_send[596] = 8'h43;
    assign to_send[597] = 8'h7a;
    assign to_send[598] = 8'h00;
    assign to_send[599] = 8'h00;
    assign to_send[600] = 8'h43;
    assign to_send[601] = 8'h53;
    assign to_send[602] = 8'h00;
    assign to_send[603] = 8'h00;
    assign to_send[604] = 8'h00;
    assign to_send[605] = 8'h00;
    assign to_send[606] = 8'h00;
    assign to_send[607] = 8'h00;
    assign to_send[608] = 8'h00;
    assign to_send[609] = 8'h00;
    assign to_send[610] = 8'h00;
    assign to_send[611] = 8'h00;
    assign to_send[612] = 8'h00;
    assign to_send[613] = 8'h00;
    assign to_send[614] = 8'h00;
    assign to_send[615] = 8'h00;
    assign to_send[616] = 8'h00;
    assign to_send[617] = 8'h00;
    assign to_send[618] = 8'h00;
    assign to_send[619] = 8'h01;
    assign to_send[620] = 8'h00;
    assign to_send[621] = 8'h00;
    assign to_send[622] = 8'h00;
    assign to_send[623] = 8'h01;
    assign to_send[624] = 8'h00;
    assign to_send[625] = 8'h00;
    assign to_send[626] = 8'h00;
    assign to_send[627] = 8'h00;
    assign to_send[628] = 8'h40;
    assign to_send[629] = 8'ha0;
    assign to_send[630] = 8'h00;
    assign to_send[631] = 8'h00;
    assign to_send[632] = 8'h41;
    assign to_send[633] = 8'h30;
    assign to_send[634] = 8'h00;
    assign to_send[635] = 8'h00;
    assign to_send[636] = 8'h42;
    assign to_send[637] = 8'h34;
    assign to_send[638] = 8'h00;
    assign to_send[639] = 8'h00;
    assign to_send[640] = 8'h00;
    assign to_send[641] = 8'h00;
    assign to_send[642] = 8'h00;
    assign to_send[643] = 8'h00;
    assign to_send[644] = 8'h42;
    assign to_send[645] = 8'h0c;
    assign to_send[646] = 8'h00;
    assign to_send[647] = 8'h00;
    assign to_send[648] = 8'h42;
    assign to_send[649] = 8'h20;
    assign to_send[650] = 8'h00;
    assign to_send[651] = 8'h00;
    assign to_send[652] = 8'h3f;
    assign to_send[653] = 8'h80;
    assign to_send[654] = 8'h00;
    assign to_send[655] = 8'h00;
    assign to_send[656] = 8'h3f;
    assign to_send[657] = 8'h80;
    assign to_send[658] = 8'h00;
    assign to_send[659] = 8'h00;
    assign to_send[660] = 8'h43;
    assign to_send[661] = 8'h7a;
    assign to_send[662] = 8'h00;
    assign to_send[663] = 8'h00;
    assign to_send[664] = 8'h43;
    assign to_send[665] = 8'h53;
    assign to_send[666] = 8'h00;
    assign to_send[667] = 8'h00;
    assign to_send[668] = 8'h43;
    assign to_send[669] = 8'h00;
    assign to_send[670] = 8'h00;
    assign to_send[671] = 8'h00;
    assign to_send[672] = 8'h00;
    assign to_send[673] = 8'h00;
    assign to_send[674] = 8'h00;
    assign to_send[675] = 8'h00;
    assign to_send[676] = 8'h00;
    assign to_send[677] = 8'h00;
    assign to_send[678] = 8'h00;
    assign to_send[679] = 8'h00;
    assign to_send[680] = 8'h00;
    assign to_send[681] = 8'h00;
    assign to_send[682] = 8'h00;
    assign to_send[683] = 8'h03;
    assign to_send[684] = 8'h00;
    assign to_send[685] = 8'h00;
    assign to_send[686] = 8'h00;
    assign to_send[687] = 8'h01;
    assign to_send[688] = 8'h00;
    assign to_send[689] = 8'h00;
    assign to_send[690] = 8'h00;
    assign to_send[691] = 8'h00;
    assign to_send[692] = 8'h41;
    assign to_send[693] = 8'hf0;
    assign to_send[694] = 8'h00;
    assign to_send[695] = 8'h00;
    assign to_send[696] = 8'h42;
    assign to_send[697] = 8'h34;
    assign to_send[698] = 8'h00;
    assign to_send[699] = 8'h00;
    assign to_send[700] = 8'h42;
    assign to_send[701] = 8'h96;
    assign to_send[702] = 8'h00;
    assign to_send[703] = 8'h00;
    assign to_send[704] = 8'h00;
    assign to_send[705] = 8'h00;
    assign to_send[706] = 8'h00;
    assign to_send[707] = 8'h00;
    assign to_send[708] = 8'h00;
    assign to_send[709] = 8'h00;
    assign to_send[710] = 8'h00;
    assign to_send[711] = 8'h00;
    assign to_send[712] = 8'h42;
    assign to_send[713] = 8'h20;
    assign to_send[714] = 8'h00;
    assign to_send[715] = 8'h00;
    assign to_send[716] = 8'h3f;
    assign to_send[717] = 8'h80;
    assign to_send[718] = 8'h00;
    assign to_send[719] = 8'h00;
    assign to_send[720] = 8'h3f;
    assign to_send[721] = 8'h80;
    assign to_send[722] = 8'h00;
    assign to_send[723] = 8'h00;
    assign to_send[724] = 8'h43;
    assign to_send[725] = 8'h7a;
    assign to_send[726] = 8'h00;
    assign to_send[727] = 8'h00;
    assign to_send[728] = 8'h43;
    assign to_send[729] = 8'h53;
    assign to_send[730] = 8'h00;
    assign to_send[731] = 8'h00;
    assign to_send[732] = 8'h43;
    assign to_send[733] = 8'h00;
    assign to_send[734] = 8'h00;
    assign to_send[735] = 8'h00;
    assign to_send[736] = 8'h00;
    assign to_send[737] = 8'h00;
    assign to_send[738] = 8'h00;
    assign to_send[739] = 8'h00;
    assign to_send[740] = 8'h00;
    assign to_send[741] = 8'h00;
    assign to_send[742] = 8'h00;
    assign to_send[743] = 8'h00;
    assign to_send[744] = 8'h00;
    assign to_send[745] = 8'h00;
    assign to_send[746] = 8'h00;
    assign to_send[747] = 8'h01;
    assign to_send[748] = 8'h00;
    assign to_send[749] = 8'h00;
    assign to_send[750] = 8'h00;
    assign to_send[751] = 8'h01;
    assign to_send[752] = 8'h00;
    assign to_send[753] = 8'h00;
    assign to_send[754] = 8'h00;
    assign to_send[755] = 8'h00;
    assign to_send[756] = 8'h41;
    assign to_send[757] = 8'hc8;
    assign to_send[758] = 8'h00;
    assign to_send[759] = 8'h00;
    assign to_send[760] = 8'h42;
    assign to_send[761] = 8'h24;
    assign to_send[762] = 8'h00;
    assign to_send[763] = 8'h00;
    assign to_send[764] = 8'h42;
    assign to_send[765] = 8'h8c;
    assign to_send[766] = 8'h00;
    assign to_send[767] = 8'h00;
    assign to_send[768] = 8'h00;
    assign to_send[769] = 8'h00;
    assign to_send[770] = 8'h00;
    assign to_send[771] = 8'h00;
    assign to_send[772] = 8'h40;
    assign to_send[773] = 8'ha0;
    assign to_send[774] = 8'h00;
    assign to_send[775] = 8'h00;
    assign to_send[776] = 8'h42;
    assign to_send[777] = 8'h20;
    assign to_send[778] = 8'h00;
    assign to_send[779] = 8'h00;
    assign to_send[780] = 8'h3f;
    assign to_send[781] = 8'h80;
    assign to_send[782] = 8'h00;
    assign to_send[783] = 8'h00;
    assign to_send[784] = 8'h3f;
    assign to_send[785] = 8'h80;
    assign to_send[786] = 8'h00;
    assign to_send[787] = 8'h00;
    assign to_send[788] = 8'h43;
    assign to_send[789] = 8'h7a;
    assign to_send[790] = 8'h00;
    assign to_send[791] = 8'h00;
    assign to_send[792] = 8'h00;
    assign to_send[793] = 8'h00;
    assign to_send[794] = 8'h00;
    assign to_send[795] = 8'h00;
    assign to_send[796] = 8'h00;
    assign to_send[797] = 8'h00;
    assign to_send[798] = 8'h00;
    assign to_send[799] = 8'h00;
    assign to_send[800] = 8'h00;
    assign to_send[801] = 8'h00;
    assign to_send[802] = 8'h00;
    assign to_send[803] = 8'h00;
    assign to_send[804] = 8'h00;
    assign to_send[805] = 8'h00;
    assign to_send[806] = 8'h00;
    assign to_send[807] = 8'h01;
    assign to_send[808] = 8'h00;
    assign to_send[809] = 8'h00;
    assign to_send[810] = 8'h00;
    assign to_send[811] = 8'h01;
    assign to_send[812] = 8'h00;
    assign to_send[813] = 8'h00;
    assign to_send[814] = 8'h00;
    assign to_send[815] = 8'h01;
    assign to_send[816] = 8'h00;
    assign to_send[817] = 8'h00;
    assign to_send[818] = 8'h00;
    assign to_send[819] = 8'h00;
    assign to_send[820] = 8'h42;
    assign to_send[821] = 8'hc8;
    assign to_send[822] = 8'h00;
    assign to_send[823] = 8'h00;
    assign to_send[824] = 8'h40;
    assign to_send[825] = 8'ha0;
    assign to_send[826] = 8'h00;
    assign to_send[827] = 8'h00;
    assign to_send[828] = 8'h43;
    assign to_send[829] = 8'h48;
    assign to_send[830] = 8'h00;
    assign to_send[831] = 8'h00;
    assign to_send[832] = 8'h00;
    assign to_send[833] = 8'h00;
    assign to_send[834] = 8'h00;
    assign to_send[835] = 8'h00;
    assign to_send[836] = 8'hc2;
    assign to_send[837] = 8'h0c;
    assign to_send[838] = 8'h00;
    assign to_send[839] = 8'h00;
    assign to_send[840] = 8'h43;
    assign to_send[841] = 8'h16;
    assign to_send[842] = 8'h00;
    assign to_send[843] = 8'h00;
    assign to_send[844] = 8'h3f;
    assign to_send[845] = 8'h80;
    assign to_send[846] = 8'h00;
    assign to_send[847] = 8'h00;
    assign to_send[848] = 8'h3f;
    assign to_send[849] = 8'h80;
    assign to_send[850] = 8'h00;
    assign to_send[851] = 8'h00;
    assign to_send[852] = 8'h43;
    assign to_send[853] = 8'h7a;
    assign to_send[854] = 8'h00;
    assign to_send[855] = 8'h00;
    assign to_send[856] = 8'h43;
    assign to_send[857] = 8'h48;
    assign to_send[858] = 8'h00;
    assign to_send[859] = 8'h00;
    assign to_send[860] = 8'h43;
    assign to_send[861] = 8'h48;
    assign to_send[862] = 8'h00;
    assign to_send[863] = 8'h00;
    assign to_send[864] = 8'h43;
    assign to_send[865] = 8'h48;
    assign to_send[866] = 8'h00;
    assign to_send[867] = 8'h00;
    assign to_send[868] = 8'h00;
    assign to_send[869] = 8'h00;
    assign to_send[870] = 8'h00;
    assign to_send[871] = 8'h00;
    assign to_send[872] = 8'h00;
    assign to_send[873] = 8'h00;
    assign to_send[874] = 8'h00;
    assign to_send[875] = 8'h03;
    assign to_send[876] = 8'h00;
    assign to_send[877] = 8'h00;
    assign to_send[878] = 8'h00;
    assign to_send[879] = 8'h01;
    assign to_send[880] = 8'h00;
    assign to_send[881] = 8'h00;
    assign to_send[882] = 8'h00;
    assign to_send[883] = 8'h00;
    assign to_send[884] = 8'h41;
    assign to_send[885] = 8'hc8;
    assign to_send[886] = 8'h00;
    assign to_send[887] = 8'h00;
    assign to_send[888] = 8'h41;
    assign to_send[889] = 8'h20;
    assign to_send[890] = 8'h00;
    assign to_send[891] = 8'h00;
    assign to_send[892] = 8'h41;
    assign to_send[893] = 8'h20;
    assign to_send[894] = 8'h00;
    assign to_send[895] = 8'h00;
    assign to_send[896] = 8'h00;
    assign to_send[897] = 8'h00;
    assign to_send[898] = 8'h00;
    assign to_send[899] = 8'h00;
    assign to_send[900] = 8'hc0;
    assign to_send[901] = 8'ha0;
    assign to_send[902] = 8'h00;
    assign to_send[903] = 8'h00;
    assign to_send[904] = 8'h00;
    assign to_send[905] = 8'h00;
    assign to_send[906] = 8'h00;
    assign to_send[907] = 8'h00;
    assign to_send[908] = 8'h3f;
    assign to_send[909] = 8'h80;
    assign to_send[910] = 8'h00;
    assign to_send[911] = 8'h00;
    assign to_send[912] = 8'h3f;
    assign to_send[913] = 8'h80;
    assign to_send[914] = 8'h00;
    assign to_send[915] = 8'h00;
    assign to_send[916] = 8'h43;
    assign to_send[917] = 8'h7a;
    assign to_send[918] = 8'h00;
    assign to_send[919] = 8'h00;
    assign to_send[920] = 8'h43;
    assign to_send[921] = 8'h53;
    assign to_send[922] = 8'h00;
    assign to_send[923] = 8'h00;
    assign to_send[924] = 8'h43;
    assign to_send[925] = 8'h00;
    assign to_send[926] = 8'h00;
    assign to_send[927] = 8'h00;
    assign to_send[928] = 8'h43;
    assign to_send[929] = 8'h00;
    assign to_send[930] = 8'h00;
    assign to_send[931] = 8'h00;
    assign to_send[932] = 8'h00;
    assign to_send[933] = 8'h00;
    assign to_send[934] = 8'h00;
    assign to_send[935] = 8'h00;
    assign to_send[936] = 8'h00;
    assign to_send[937] = 8'h00;
    assign to_send[938] = 8'h00;
    assign to_send[939] = 8'h03;
    assign to_send[940] = 8'h00;
    assign to_send[941] = 8'h00;
    assign to_send[942] = 8'h00;
    assign to_send[943] = 8'h02;
    assign to_send[944] = 8'h00;
    assign to_send[945] = 8'h00;
    assign to_send[946] = 8'h00;
    assign to_send[947] = 8'h00;
    assign to_send[948] = 8'h41;
    assign to_send[949] = 8'hc8;
    assign to_send[950] = 8'h00;
    assign to_send[951] = 8'h00;
    assign to_send[952] = 8'h41;
    assign to_send[953] = 8'ha0;
    assign to_send[954] = 8'h00;
    assign to_send[955] = 8'h00;
    assign to_send[956] = 8'h41;
    assign to_send[957] = 8'ha0;
    assign to_send[958] = 8'h00;
    assign to_send[959] = 8'h00;
    assign to_send[960] = 8'h00;
    assign to_send[961] = 8'h00;
    assign to_send[962] = 8'h00;
    assign to_send[963] = 8'h00;
    assign to_send[964] = 8'h00;
    assign to_send[965] = 8'h00;
    assign to_send[966] = 8'h00;
    assign to_send[967] = 8'h00;
    assign to_send[968] = 8'h42;
    assign to_send[969] = 8'h8c;
    assign to_send[970] = 8'h00;
    assign to_send[971] = 8'h00;
    assign to_send[972] = 8'h3f;
    assign to_send[973] = 8'h80;
    assign to_send[974] = 8'h00;
    assign to_send[975] = 8'h00;
    assign to_send[976] = 8'h3e;
    assign to_send[977] = 8'h99;
    assign to_send[978] = 8'h99;
    assign to_send[979] = 8'h9a;
    assign to_send[980] = 8'h00;
    assign to_send[981] = 8'h00;
    assign to_send[982] = 8'h00;
    assign to_send[983] = 8'h00;
    assign to_send[984] = 8'h00;
    assign to_send[985] = 8'h00;
    assign to_send[986] = 8'h00;
    assign to_send[987] = 8'h00;
    assign to_send[988] = 8'h00;
    assign to_send[989] = 8'h00;
    assign to_send[990] = 8'h00;
    assign to_send[991] = 8'h00;
    assign to_send[992] = 8'h43;
    assign to_send[993] = 8'h7f;
    assign to_send[994] = 8'h00;
    assign to_send[995] = 8'h00;
    assign to_send[996] = 8'h00;
    assign to_send[997] = 8'h00;
    assign to_send[998] = 8'h00;
    assign to_send[999] = 8'h02;
    assign to_send[1000] = 8'h00;
    assign to_send[1001] = 8'h00;
    assign to_send[1002] = 8'h00;
    assign to_send[1003] = 8'h03;
    assign to_send[1004] = 8'h00;
    assign to_send[1005] = 8'h00;
    assign to_send[1006] = 8'h00;
    assign to_send[1007] = 8'h01;
    assign to_send[1008] = 8'h00;
    assign to_send[1009] = 8'h00;
    assign to_send[1010] = 8'h00;
    assign to_send[1011] = 8'h00;
    assign to_send[1012] = 8'h41;
    assign to_send[1013] = 8'ha0;
    assign to_send[1014] = 8'h00;
    assign to_send[1015] = 8'h00;
    assign to_send[1016] = 8'h41;
    assign to_send[1017] = 8'ha0;
    assign to_send[1018] = 8'h00;
    assign to_send[1019] = 8'h00;
    assign to_send[1020] = 8'h41;
    assign to_send[1021] = 8'ha0;
    assign to_send[1022] = 8'h00;
    assign to_send[1023] = 8'h00;
    assign to_send[1024] = 8'h42;
    assign to_send[1025] = 8'hc8;
    assign to_send[1026] = 8'h00;
    assign to_send[1027] = 8'h00;
    assign to_send[1028] = 8'h42;
    assign to_send[1029] = 8'h20;
    assign to_send[1030] = 8'h00;
    assign to_send[1031] = 8'h00;
    assign to_send[1032] = 8'h42;
    assign to_send[1033] = 8'hf0;
    assign to_send[1034] = 8'h00;
    assign to_send[1035] = 8'h00;
    assign to_send[1036] = 8'h3f;
    assign to_send[1037] = 8'h80;
    assign to_send[1038] = 8'h00;
    assign to_send[1039] = 8'h00;
    assign to_send[1040] = 8'h3f;
    assign to_send[1041] = 8'h80;
    assign to_send[1042] = 8'h00;
    assign to_send[1043] = 8'h00;
    assign to_send[1044] = 8'h43;
    assign to_send[1045] = 8'h16;
    assign to_send[1046] = 8'h00;
    assign to_send[1047] = 8'h00;
    assign to_send[1048] = 8'h43;
    assign to_send[1049] = 8'h7f;
    assign to_send[1050] = 8'h00;
    assign to_send[1051] = 8'h00;
    assign to_send[1052] = 8'h43;
    assign to_send[1053] = 8'h7f;
    assign to_send[1054] = 8'h00;
    assign to_send[1055] = 8'h00;
    assign to_send[1056] = 8'h43;
    assign to_send[1057] = 8'h7f;
    assign to_send[1058] = 8'h00;
    assign to_send[1059] = 8'h00;
    assign to_send[1060] = 8'h00;
    assign to_send[1061] = 8'h00;
    assign to_send[1062] = 8'h00;
    assign to_send[1063] = 8'h00;
    assign to_send[1064] = 8'h00;
    assign to_send[1065] = 8'h00;
    assign to_send[1066] = 8'h00;
    assign to_send[1067] = 8'h02;
    assign to_send[1068] = 8'h00;
    assign to_send[1069] = 8'h00;
    assign to_send[1070] = 8'h00;
    assign to_send[1071] = 8'h02;
    assign to_send[1072] = 8'h00;
    assign to_send[1073] = 8'h00;
    assign to_send[1074] = 8'h00;
    assign to_send[1075] = 8'h00;
    assign to_send[1076] = 8'h00;
    assign to_send[1077] = 8'h00;
    assign to_send[1078] = 8'h00;
    assign to_send[1079] = 8'h00;
    assign to_send[1080] = 8'h00;
    assign to_send[1081] = 8'h00;
    assign to_send[1082] = 8'h00;
    assign to_send[1083] = 8'h00;
    assign to_send[1084] = 8'hbf;
    assign to_send[1085] = 8'h80;
    assign to_send[1086] = 8'h00;
    assign to_send[1087] = 8'h00;
    assign to_send[1088] = 8'h00;
    assign to_send[1089] = 8'h00;
    assign to_send[1090] = 8'h00;
    assign to_send[1091] = 8'h00;
    assign to_send[1092] = 8'h00;
    assign to_send[1093] = 8'h00;
    assign to_send[1094] = 8'h00;
    assign to_send[1095] = 8'h00;
    assign to_send[1096] = 8'h43;
    assign to_send[1097] = 8'h48;
    assign to_send[1098] = 8'h00;
    assign to_send[1099] = 8'h00;
    assign to_send[1100] = 8'h3f;
    assign to_send[1101] = 8'h80;
    assign to_send[1102] = 8'h00;
    assign to_send[1103] = 8'h00;
    assign to_send[1104] = 8'h3e;
    assign to_send[1105] = 8'h4c;
    assign to_send[1106] = 8'hcc;
    assign to_send[1107] = 8'hcd;
    assign to_send[1108] = 8'h00;
    assign to_send[1109] = 8'h00;
    assign to_send[1110] = 8'h00;
    assign to_send[1111] = 8'h00;
    assign to_send[1112] = 8'h43;
    assign to_send[1113] = 8'h7f;
    assign to_send[1114] = 8'h00;
    assign to_send[1115] = 8'h00;
    assign to_send[1116] = 8'h00;
    assign to_send[1117] = 8'h00;
    assign to_send[1118] = 8'h00;
    assign to_send[1119] = 8'h00;
    assign to_send[1120] = 8'h00;
    assign to_send[1121] = 8'h00;
    assign to_send[1122] = 8'h00;
    assign to_send[1123] = 8'h00;
    assign to_send[1124] = 8'hff;
    assign to_send[1125] = 8'hff;
    assign to_send[1126] = 8'hff;
    assign to_send[1127] = 8'hff;
    assign to_send[1128] = 8'h00;
    assign to_send[1129] = 8'h00;
    assign to_send[1130] = 8'h00;
    assign to_send[1131] = 8'h00;
    assign to_send[1132] = 8'h00;
    assign to_send[1133] = 8'h00;
    assign to_send[1134] = 8'h00;
    assign to_send[1135] = 8'h01;
    assign to_send[1136] = 8'h00;
    assign to_send[1137] = 8'h00;
    assign to_send[1138] = 8'h00;
    assign to_send[1139] = 8'h02;
    assign to_send[1140] = 8'hff;
    assign to_send[1141] = 8'hff;
    assign to_send[1142] = 8'hff;
    assign to_send[1143] = 8'hff;
    assign to_send[1144] = 8'h00;
    assign to_send[1145] = 8'h00;
    assign to_send[1146] = 8'h00;
    assign to_send[1147] = 8'h03;
    assign to_send[1148] = 8'h00;
    assign to_send[1149] = 8'h00;
    assign to_send[1150] = 8'h00;
    assign to_send[1151] = 8'h01;
    assign to_send[1152] = 8'h00;
    assign to_send[1153] = 8'h00;
    assign to_send[1154] = 8'h00;
    assign to_send[1155] = 8'h04;
    assign to_send[1156] = 8'hff;
    assign to_send[1157] = 8'hff;
    assign to_send[1158] = 8'hff;
    assign to_send[1159] = 8'hff;
    assign to_send[1160] = 8'h00;
    assign to_send[1161] = 8'h00;
    assign to_send[1162] = 8'h00;
    assign to_send[1163] = 8'h05;
    assign to_send[1164] = 8'h00;
    assign to_send[1165] = 8'h00;
    assign to_send[1166] = 8'h00;
    assign to_send[1167] = 8'h06;
    assign to_send[1168] = 8'h00;
    assign to_send[1169] = 8'h00;
    assign to_send[1170] = 8'h00;
    assign to_send[1171] = 8'h07;
    assign to_send[1172] = 8'hff;
    assign to_send[1173] = 8'hff;
    assign to_send[1174] = 8'hff;
    assign to_send[1175] = 8'hff;
    assign to_send[1176] = 8'h00;
    assign to_send[1177] = 8'h00;
    assign to_send[1178] = 8'h00;
    assign to_send[1179] = 8'h08;
    assign to_send[1180] = 8'hff;
    assign to_send[1181] = 8'hff;
    assign to_send[1182] = 8'hff;
    assign to_send[1183] = 8'hff;
    assign to_send[1184] = 8'h00;
    assign to_send[1185] = 8'h00;
    assign to_send[1186] = 8'h00;
    assign to_send[1187] = 8'h09;
    assign to_send[1188] = 8'h00;
    assign to_send[1189] = 8'h00;
    assign to_send[1190] = 8'h00;
    assign to_send[1191] = 8'h0a;
    assign to_send[1192] = 8'hff;
    assign to_send[1193] = 8'hff;
    assign to_send[1194] = 8'hff;
    assign to_send[1195] = 8'hff;
    assign to_send[1196] = 8'h00;
    assign to_send[1197] = 8'h00;
    assign to_send[1198] = 8'h00;
    assign to_send[1199] = 8'h0c;
    assign to_send[1200] = 8'hff;
    assign to_send[1201] = 8'hff;
    assign to_send[1202] = 8'hff;
    assign to_send[1203] = 8'hff;
    assign to_send[1204] = 8'h00;
    assign to_send[1205] = 8'h00;
    assign to_send[1206] = 8'h00;
    assign to_send[1207] = 8'h0d;
    assign to_send[1208] = 8'hff;
    assign to_send[1209] = 8'hff;
    assign to_send[1210] = 8'hff;
    assign to_send[1211] = 8'hff;
    assign to_send[1212] = 8'h00;
    assign to_send[1213] = 8'h00;
    assign to_send[1214] = 8'h00;
    assign to_send[1215] = 8'h0e;
    assign to_send[1216] = 8'hff;
    assign to_send[1217] = 8'hff;
    assign to_send[1218] = 8'hff;
    assign to_send[1219] = 8'hff;
    assign to_send[1220] = 8'h00;
    assign to_send[1221] = 8'h00;
    assign to_send[1222] = 8'h00;
    assign to_send[1223] = 8'h0f;
    assign to_send[1224] = 8'hff;
    assign to_send[1225] = 8'hff;
    assign to_send[1226] = 8'hff;
    assign to_send[1227] = 8'hff;
    assign to_send[1228] = 8'h00;
    assign to_send[1229] = 8'h00;
    assign to_send[1230] = 8'h00;
    assign to_send[1231] = 8'h10;
    assign to_send[1232] = 8'hff;
    assign to_send[1233] = 8'hff;
    assign to_send[1234] = 8'hff;
    assign to_send[1235] = 8'hff;
    assign to_send[1236] = 8'hff;
    assign to_send[1237] = 8'hff;
    assign to_send[1238] = 8'hff;
    assign to_send[1239] = 8'hff;
    assign to_send[1240] = 8'h00;
    assign to_send[1241] = 8'h00;
    assign to_send[1242] = 8'h00;
    assign to_send[1243] = 8'h0b;
    assign to_send[1244] = 8'h00;
    assign to_send[1245] = 8'h00;
    assign to_send[1246] = 8'h00;
    assign to_send[1247] = 8'h00;
    assign to_send[1248] = 8'h00;
    assign to_send[1249] = 8'h00;
    assign to_send[1250] = 8'h00;
    assign to_send[1251] = 8'h01;
    assign to_send[1252] = 8'h00;
    assign to_send[1253] = 8'h00;
    assign to_send[1254] = 8'h00;
    assign to_send[1255] = 8'h02;
    assign to_send[1256] = 8'h00;
    assign to_send[1257] = 8'h00;
    assign to_send[1258] = 8'h00;
    assign to_send[1259] = 8'h03;
    assign to_send[1260] = 8'h00;
    assign to_send[1261] = 8'h00;
    assign to_send[1262] = 8'h00;
    assign to_send[1263] = 8'h04;
    assign to_send[1264] = 8'h00;
    assign to_send[1265] = 8'h00;
    assign to_send[1266] = 8'h00;
    assign to_send[1267] = 8'h06;
    assign to_send[1268] = 8'hff;
    assign to_send[1269] = 8'hff;
    assign to_send[1270] = 8'hff;
    assign to_send[1271] = 8'hff;
    assign to_send[1272] = 8'h00;
    assign to_send[1273] = 8'h00;
    assign to_send[1274] = 8'h00;
    assign to_send[1275] = 8'h63;
    assign to_send[1276] = 8'h00;
    assign to_send[1277] = 8'h00;
    assign to_send[1278] = 8'h00;
    assign to_send[1279] = 8'h09;
    assign to_send[1280] = 8'h00;
    assign to_send[1281] = 8'h00;
    assign to_send[1282] = 8'h00;
    assign to_send[1283] = 8'h08;
    assign to_send[1284] = 8'h00;
    assign to_send[1285] = 8'h00;
    assign to_send[1286] = 8'h00;
    assign to_send[1287] = 8'h07;
    assign to_send[1288] = 8'h00;
    assign to_send[1289] = 8'h00;
    assign to_send[1290] = 8'h00;
    assign to_send[1291] = 8'h05;
    assign to_send[1292] = 8'hff;
    assign to_send[1293] = 8'hff;
    assign to_send[1294] = 8'hff;
    assign to_send[1295] = 8'hff;
    assign to_send[1296] = 8'hff;
    assign to_send[1297] = 8'hff;
    assign to_send[1298] = 8'hff;
    assign to_send[1299] = 8'hff;

    reg [32-1:0] idx;
    reg started;
    reg order;
    wire sendable;

    always @(posedge clk) begin
        if (~rstn) begin
            order <= 1'b0;
            started <= 1'b0;
            idx <=32'b0;
        end else if (sendable) begin
            if (started && (idx<32'd1300)) begin
                idx <= idx + 32'b1;
            end else begin
                started <= 1'b1;
            end
            if (idx<32'd1300) begin
                order <= 1'b1;
            end else begin
                order <= 1'b0;
            end
        end else begin
            order <= 1'b0;
        end
    end

    uart_tx #(CLK_FREQ, BAUD)
    m_uart_tx(
        order, to_send[idx], sendable, rx, clk, rstn);

endmodule

`default_nettype wire
